*FD

.include spice_lib/sky130.lib

xm1 1 2 3 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm2 0 2 3 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm3 3 clkb 4 1 sky130_fd_pr__pfet_01v8 l=150n w=420n
xm4 3 clk 4 0 sky130_fd_pr__nfet_01v8 l=150n w=840n

xm7 1 4 5 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm8 0 4 5 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm9 5 clk 6 1 sky130_fd_pr__pfet_01v8 l=150n w=420n
xm10 5 clkb 6 0 sky130_fd_pr__nfet_01v8 l=150n w=640n

xm11 1 6 2 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm12 0 6 2 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm13 1 clk clkb 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm14 0 clk clkb 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

v1 1 0 1.8
v2 clk 0 PULSE 0 1.8 1n 6p 6p 5ns 10ns

c1 6 0 10f
.control
tran 0.1ns 0.2us
plot v(6) v(clk)+2
.endc

.end

